`timescale 1ns/1ps
module cu(
    input rst,
    input branch_predict_success,
    input branch_predict_fail,
    input [31:0] rf_rdata1,
    input [31:0] rf_rdata2,
    input [4:0] rs,
    input [4:0] rt,
    input [4:0] rd,
    input [4:0] shamt,
    input [15:0] immediate,
    input [25:0] address,
    input [7:0] INST,
    input [31:0] pc4,
    input [31:0] ext18,
    input [31:0] cp0_exec_addr,
    input [5:0] cp0_int_i, 
    input [31:0] cp0_status,
    input LLbit_odata,
    output reg DMEM_wena,
    output reg [3:0] data_type,
    output reg CBW_sign,
    output reg CHW_sign,
    output reg [7:0] mux_pc,
    output reg [7:0] mux_rf,
    output reg mux_rf_DMEM,
    output reg [7:0] mux_alu,
    output reg [7:0] mux_hi,
    output reg [7:0] mux_lo,
    output reg rf_wena,
    output reg [3:0] mov_cond,
    output reg [4:0] rf_waddr,
    output reg [3:0] alu_aluc,
    output reg hi_ena,
    output reg lo_ena,
    output reg [3:0] hi_lo_func,
    output reg EXT1_n_c,
    output reg EXT16_sign,
    output mfc0,
    output mtc0,
    output reg exception,
    output eret,
    output reg [4:0] cause,
    output reg blockade,
    output branch_inst,
    output branch_predict,
    output reg [3:0] branch_flag,
    output reg [31:0] branch_fail_pc,
    output reg LLbit_idata,
    output reg LLbit_wena
);
    wire [31:0] ext16;
    //assign branch_predict=0;
    predictor PREDICTOR(
        .rst(rst),
        .success(branch_predict_success),
        .fail(branch_predict_fail),
        .branch_predict(branch_predict)
    );
    parameter Wdata=4'd0,Hdata=4'd1,Bdata=4'd2,Ldata=4'd3,Rdata=4'd4;
    parameter ADD=8'd1,ADDU=8'd2,SUB=8'd3,SUBU=8'd4,AND=8'd5,OR=8'd6,XOR=8'd7,NOR=8'd8,SLT=8'd9,SLTU=8'd10,SLL=8'd11,SRL=8'd12,SRA=8'd13,SLLV=8'd14,SRLV=8'd15,SRAV=8'd16,JR=8'd17,
    ADDI=8'd18,ADDIU=8'd19,ANDI=8'd20,ORI=8'd21,XORI=8'd22,LW=8'd23,SW=8'd24,BEQ=8'd25,BNE=8'd26,SLTI=8'd27,SLTIU=8'd28,LUI=8'd29,J=8'd30,JAL=8'd31,
    DIV=8'd32,DIVU=8'd33,MULT=8'd34,MULTU=8'd35,BGEZ=8'd36,JALR=8'd37,LBU=8'd38,LHU=8'd39,LB=8'd40,LH=8'd41,SB=8'd42,SH=8'd43,BREAK=8'd44,SYSCALL=8'd45,ERET=8'd46,MFHI=8'd47,MFLO=8'd48,
    MTHI=8'd49,MTLO=8'd50,MFC0=8'd51,MTC0=8'd52,CLZ=8'd53,TEQ=8'd54,MUL=8'd55,
    MOVN=8'd56,MOVZ=8'd57,CLO=8'd58,MADD=8'd59,MADDU=8'd60,MSUB=8'd61,MSUBU=8'd62,BGEZAL=8'd63,BGTZ=8'd64,BLEZ=8'd65,BLTZ=8'd66,BLTZAL=8'd67,
    LL=8'd68,LWL=8'd69,LWR=8'd70,SC=8'd71,SWL=8'd72,SWR=8'd73,TGE=8'd74,TGEU=8'd75,TLT=8'd76,TLTU=8'd77,TNE=8'd78,TEQI=8'd79,TGEI=8'd80,TGEIU=8'd81,TLTI=8'd82,TLTIU=8'd83,TNEI=8'd84;
    parameter mux_pc_NPC=8'd0,mux_pc_Rs=8'd1,mux_pc_EXT18=8'd2,mux_pc_II=8'd3,mux_pc_EPC=8'd4;
    parameter mux_rf_ALU=8'd0,mux_rf_EXT1=8'd1,mux_rf_PC=8'd2,mux_rf_CLZ=8'd3,mux_rf_HI=8'd4,mux_rf_LO=8'd5,mux_rf_CPR=8'd6,mux_rf_MUL=8'd7,mux_rf_CLO=8'd8,mux_rf_O=8'd9,mux_rf_Z=8'd10;
    parameter mux_alu_Rs_Rt=8'd0,mux_alu_ext5_Rt=8'd1,mux_alu_Rs_EXT16=8'd2,mux_alu_x_EXT16=8'd3,mux_alu_Rs_0=8'd4;
    parameter mux_hi_Rs=8'd0,mux_hi_DIV=8'd1,mux_hi_DIVU=8'd2,mux_hi_MULT=8'd3,mux_hi_MULTU=8'd4;
    parameter mux_lo_Rs=8'd0,mux_lo_DIV=8'd1,mux_lo_DIVU=8'd2,mux_lo_MULT=8'd3,mux_lo_MULTU=8'd4;
    parameter EXC_Int=5'd0,EXC_Sys=5'd8,EXC_Bp=5'd9,EXC_RI=5'd10,EXC_Ov=5'd12,EXC_Tr=5'd13;//EXC_syscall=5'b01000,EXC_break=5'b01001,EXC_teq=5'b01101;
    parameter branch_NONE=4'd0,branch_BEQ=4'd1,branch_BNE=4'd2,branch_BGEZ=4'd3,
    branch_BGTZ=4'd5,branch_BLEZ=4'd6,branch_BLTZ=4'd7;
    parameter mov_cond_NONE=4'd0,mov_cond_N=4'd1,mov_cond_Z=4'd2;
    parameter hi_lo_func_NONE=4'd0,hi_lo_func_MADD=4'd1,hi_lo_func_MADDU=4'd2,hi_lo_func_MSUB=4'd3,hi_lo_func_MSUBU=4'd4;
    assign mfc0=(INST==MFC0);
    assign mtc0=(INST==MTC0);
    //assign exception=(cp0_int_i!=6'd0)|(INST==BREAK)|(INST==SYSCALL)|(INST==ERET)|(INST==TEQ)|(INST>=TGE&&INST<=TNEI);
    assign eret=(INST==ERET);
    assign branch_inst=(INST==BEQ)|(INST==BNE)|(INST==BGEZ)|(INST>=BGEZAL&&INST<=BLTZAL);
    assign ext16={{16{immediate[15]}},immediate};
    always@(*)
    begin
        //if(cp0_int_i[0]&&cp0_status[0]&~cp0_status[1]&cp0_status[10])//timer_int
        if(cp0_int_i[0])
        begin
            exception<=1;
            DMEM_wena<=0;
            data_type<=4'bx; 
            CBW_sign<=1'bx;
            CHW_sign<=1'bx; 
            mux_pc<=mux_pc_EPC;
            mux_rf<=8'bx;
            mux_rf_DMEM<=1'bx;
            mux_alu<=8'bx;
            mux_hi<=8'bx;
            mux_lo<=8'bx;
            rf_wena<=0;
            mov_cond<=mov_cond_NONE;
            rf_waddr<=5'bx;
            alu_aluc<=4'bx;
            hi_ena<=0;
            lo_ena<=0;
            hi_lo_func<=hi_lo_func_NONE;
            EXT1_n_c<=1'bx;
            EXT16_sign<=1'bx;
            cause<=EXC_Int;
            blockade<=1;
            branch_flag<=branch_NONE;
            branch_fail_pc<=32'bx;
            LLbit_idata<=1'bx;
            LLbit_wena<=0;
        end
        else
        begin
        case(INST)
            //#1
            ADD:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx;
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;            
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#2
            ADDU:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0000;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#3
            SUB:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0011;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#4
            SUBU:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0001;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#5
            AND:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0100;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#6
            OR:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0101;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#7
            XOR:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0110;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#8
            NOR:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b0111;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#9
            SLT:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_EXT1;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1011;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=0;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#10
            SLTU:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_EXT1;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#11
            SLL:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx;
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;  
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_ext5_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b111x;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#12
            SRL:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_ext5_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1101;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#13
            SRA:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_ext5_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1100;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#14
            SLLV:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b111x;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#15
            SRLV:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1101;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#16
            SRAV:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_Rt;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'b1100;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#17
            JR:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_Rs;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#18
            ADDI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#19
            ADDIU:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0000;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#20
            ANDI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0100;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=0;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#21
            ORI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0101;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=0;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#22
            XORI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0110;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=0;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#23
            LW:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=Wdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#24
            SW:begin
                exception<=0;
                DMEM_wena<=1;
                data_type<=Wdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#25
            BEQ:begin
                exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BEQ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BEQ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#26
            BNE:begin
                exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BNE;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BNE;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#27
            SLTI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_EXT1;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b1011;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=0;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#28
            SLTIU:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_EXT1;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b1010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1;
                EXT16_sign<=0;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#29
            LUI:begin
                exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_x_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b100x;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=0;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#30
            J:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_II;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#31
            JAL:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx;
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;  
                mux_pc<=mux_pc_II;
                mux_rf<=mux_rf_PC;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'd31;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#32
            DIV:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_DIV;
                mux_lo<=mux_lo_DIV;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#33
            DIVU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_DIVU;
                mux_lo<=mux_lo_DIVU;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#34
            MULT:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULT;
                mux_lo<=mux_lo_MULT;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#35
            MULTU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULTU;
                mux_lo<=mux_lo_MULTU;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#36
            BGEZ:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BGEZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BGEZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end        
            //#37
            JALR:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_Rs;
                mux_rf<=mux_rf_PC;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#38
            LBU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Bdata; 
                CBW_sign<=0;
                CHW_sign<=0; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#39
            LHU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Hdata; 
                CBW_sign<=0;
                CHW_sign<=0;
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#40
            LB:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Bdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#41
            LH:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Hdata; 
                CBW_sign<=1;
                CHW_sign<=1;
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#42
            SB:begin
				exception<=0;
                DMEM_wena<=1;
                data_type<=Bdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#43
            SH:begin
				exception<=0;
                DMEM_wena<=1;
                data_type<=Hdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#44
            BREAK:begin
                exception<=1;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_EPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=EXC_Bp;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#45
            SYSCALL:begin
                exception<=1;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_EPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=EXC_Sys;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //$46
            ERET:begin
                exception<=1;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_EPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=1;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#47
            MFHI:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_HI;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#48
            MFLO:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_LO;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#49
            MTHI:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_Rs;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#50
            MTLO:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=mux_lo_Rs;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#51
            MFC0:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_CPR;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#52
            MTC0:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#53
            CLZ:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_CLZ;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#54
            TEQ:begin
                if(rf_rdata1==rf_rdata2)
                begin
                    exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#55
            MUL:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_MUL;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#56
            MOVN:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx;
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;            
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_0;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_N;
                rf_waddr<=rd;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#57
            MOVZ:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx;
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;            
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_ALU;
                mux_rf_DMEM<=0;
                mux_alu<=mux_alu_Rs_0;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_Z;
                rf_waddr<=rd;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#58
            CLO:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx;
                mux_pc<=mux_pc_NPC;
                mux_rf<=mux_rf_CLO;
                mux_rf_DMEM<=0;
                mux_alu<=8'bx;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rd;
                alu_aluc<=4'bx;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#59
            MADD:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULT;
                mux_lo<=mux_lo_MULT;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_MADD;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#60
            MADDU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULTU;
                mux_lo<=mux_lo_MULTU;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_MADDU;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#61
            MSUB:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULT;
                mux_lo<=mux_lo_MULT;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_MSUB;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#62
            MSUBU:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=4'bx; 
                CBW_sign<=1'bx;
                CHW_sign<=1'bx; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=8'bx;
                mux_hi<=mux_hi_MULTU;
                mux_lo<=mux_lo_MULTU;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'bx;
                hi_ena<=1;
                lo_ena<=1;
                hi_lo_func<=hi_lo_func_MSUBU;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1'bx;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#63
            BGTZ:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BGTZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BGTZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#64
            BLEZ:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BLEZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BLEZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#65
            BLTZ:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BLTZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BLTZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#66
            BLTZAL:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=mux_rf_PC;
                    mux_rf_DMEM<=0;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'd31;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BLTZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=mux_rf_PC;
                    mux_rf_DMEM<=0;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'd31;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BLTZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#67
            BGEZAL:begin
				exception<=0;
                if(branch_predict)
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_EXT18;
                    mux_rf<=mux_rf_PC;
                    mux_rf_DMEM<=0;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'd31;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=1;
                    branch_flag<=branch_BGEZ;
                    branch_fail_pc<=pc4;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=mux_rf_PC;
                    mux_rf_DMEM<=0;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'd31;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_BGEZ;
                    branch_fail_pc<=ext18;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#68
            LWL:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Ldata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end 
            //#69
            LWR:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Rdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end      
            //#70
            SWL:begin
				exception<=0;
                DMEM_wena<=1;
                data_type<=Ldata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end 
            //#71
            SWR:begin
				exception<=0;
                DMEM_wena<=1;
                data_type<=Rdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1'bx;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=0;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=5'bx;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'bx;
                LLbit_wena<=0;
            end
            //#72
            LL:begin
				exception<=0;
                DMEM_wena<=0;
                data_type<=Wdata; 
                CBW_sign<=1;
                CHW_sign<=1; 
                mux_pc<=mux_pc_NPC;
                mux_rf<=8'bx;
                mux_rf_DMEM<=1;
                mux_alu<=mux_alu_Rs_EXT16;
                mux_hi<=8'bx;
                mux_lo<=8'bx;
                rf_wena<=1;
                mov_cond<=mov_cond_NONE;
                rf_waddr<=rt;
                alu_aluc<=4'b0010;
                hi_ena<=0;
                lo_ena<=0;
                hi_lo_func<=hi_lo_func_NONE;
                EXT1_n_c<=1'bx;
                EXT16_sign<=1;
                cause<=5'bx;
                blockade<=0;
                branch_flag<=branch_NONE;
                branch_fail_pc<=32'bx;
                LLbit_idata<=1'b1;
                LLbit_wena<=1;
            end
            //#73
            SC:begin
				exception<=0;
                if(LLbit_odata)
                begin
                    DMEM_wena<=1;
                    data_type<=Wdata;
                    CBW_sign<=1;
                    CHW_sign<=1; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=mux_rf_O;
                    mux_rf_DMEM<=0;
                    mux_alu<=mux_alu_Rs_EXT16;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=rt;
                    alu_aluc<=4'b0010;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
                    DMEM_wena<=0;
                    data_type<=4'bx;
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx; 
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=mux_rf_Z;
                    mux_rf_DMEM<=0;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=1;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=rt;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=5'bx;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#74
            TGE:begin
                if((rf_rdata1[31]==rf_rdata2[31]&&rf_rdata1>=rf_rdata2)||(rf_rdata1[31]==0&&rf_rdata2[31]==1))
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#75
            TGEU:begin
                if(rf_rdata1>=rf_rdata2)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#76
            TLT:begin
                if((rf_rdata1[31]==rf_rdata2[31]&&rf_rdata1<rf_rdata2)||(rf_rdata1[31]==1&&rf_rdata2[31]==0))
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#77
            TLTU:begin
                if(rf_rdata1<rf_rdata2)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#78
            TNE:begin
                if(rf_rdata1!=rf_rdata2)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#79
            TEQI:begin
                if(rf_rdata1==ext16)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#80
            TGEI:begin
                if((rf_rdata1[31]==ext16[31]&&rf_rdata1>=ext16)||(rf_rdata1[31]==0&&ext16[31]==1))
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#81
            TGEIU:begin
                if(rf_rdata1>=ext16)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#82
            TLTI:begin
                if((rf_rdata1[31]==ext16[31]&&rf_rdata1<ext16)||(rf_rdata1[31]==1&&ext16[31]==0))
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#83
            TLTIU:begin
                if(rf_rdata1<ext16)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
            //#84
            TNEI:begin
                if(rf_rdata1!=ext16)
                begin
					exception<=1;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;
                    mux_pc<=mux_pc_EPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=1;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
                else
                begin
					exception<=0;
                    DMEM_wena<=0;
                    data_type<=4'bx; 
                    CBW_sign<=1'bx;
                    CHW_sign<=1'bx;                     
                    mux_pc<=mux_pc_NPC;
                    mux_rf<=8'bx;
                    mux_rf_DMEM<=1'bx;
                    mux_alu<=8'bx;
                    mux_hi<=8'bx;
                    mux_lo<=8'bx;
                    rf_wena<=0;
                    mov_cond<=mov_cond_NONE;
                    rf_waddr<=5'bx;
                    alu_aluc<=4'bx;
                    hi_ena<=0;
                    lo_ena<=0;
                    hi_lo_func<=hi_lo_func_NONE;
                    EXT1_n_c<=1'bx;
                    EXT16_sign<=1'bx;
                    cause<=EXC_Tr;
                    blockade<=0;
                    branch_flag<=branch_NONE;
                    branch_fail_pc<=32'bx;
                    LLbit_idata<=1'bx;
                    LLbit_wena<=0;
                end
            end
        endcase
        end
    end
endmodule